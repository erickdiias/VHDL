--
--
--
--

library ieee;
use ieee.std_logic_1164.all;

entity HCRS04 is
    port();
end entity;

architecture main of HCRS04 is
begin
end architecture;