entity semaforos 